V1 0 1 dc 15
R1 2 3 0.068181
R2 4 5 0.089932
R3 6 7 0.087560
R4 8 9 0.043529
R5 10 11 0.064742
R6 12 13 0.044420
R7 14 15 0.071837
R8 16 17 0.184061
R9 18 1 0.064941
R10 19 20 0.071267
R11 21 22 0.075622
R12 23 1 0.064672
R13 24 25 0.055011
R14 0 26 0.061432
R15 27 28 0.068416
R16 29 30 0.079033
R17 31 32 0.149925
R18 0 33 0.106829
R19 9 2 0.029860
R20 3 14 0.015013
R21 3 19 0.100575
R22 5 19 0.017832
R23 26 4 0.039886
R24 33 4 0.013583
R25 17 6 0.011612
R26 9 24 0.013808
R27 9 27 0.024336
R28 15 10 0.009895
R29 11 18 0.031260
R30 13 16 0.034322
R31 28 12 0.028444
R32 25 14 0.024463
R33 28 14 0.016237
R34 17 18 0.044077
R35 25 16 0.081811
R36 28 16 0.036152
R37 20 21 0.048043
R38 20 23 0.007903
R39 30 19 0.023751
R40 26 29 0.015652
R41 32 27 0.014558
.dc V1 15 15 1
.print dc i(V1)
.end
