V1 0 1 dc 15
R1 2 3 0.055139
R2 4 1 0.059797
R3 0 5 0.080647
R4 6 7 0.064689
R5 8 9 0.118648
R6 0 10 0.188375
R7 11 12 0.096978
R8 0 13 0.084129
R9 14 15 0.079598
R10 16 1 0.090438
R11 17 18 0.078540
R12 19 1 0.101922
R13 20 21 0.042327
R14 22 23 0.106572
R15 0 24 0.045727
R16 25 26 0.054545
R17 0 27 0.084956
R18 28 1 0.075453
R19 7 2 0.026965
R20 3 16 0.091951
R21 21 2 0.030288
R22 3 22 0.023197
R23 3 25 0.012738
R24 26 4 0.013944
R25 5 14 0.017123
R26 7 22 0.037138
R27 27 6 0.010751
R28 13 8 0.022347
R29 9 16 0.037333
R30 9 17 0.023946
R31 10 11 0.036182
R32 10 20 0.038995
R33 13 11 0.013647
R34 12 16 0.012154
R35 15 17 0.029365
R36 18 19 0.016349
R37 24 20 0.006650
R38 23 28 0.015265
.dc V1 15 15 1
.print dc i(V1)
.end
